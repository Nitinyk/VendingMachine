`include "transaction.sv"
`include "generator.sv"
`include "cov.sv"
`include "bfm.sv"
`include "interface.sv"
`include "environment.sv"
`include "test.sv"
`include "design.sv"
`include "testbench_top.sv"
`include "monitor.sv"
//`include "scoreboard.sv"
