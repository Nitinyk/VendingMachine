`include "environment.sv"
`include "scoreboard.sv"
`include "transaction.sv"
`include "generator.sv"
`include "interface.sv"
`include "test.sv"
`include "design.sv"
`include "tb_top.sv"
`include "driver.sv"
`include "monitor.sv"
