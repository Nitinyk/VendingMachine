 class transaction;

//only input signals for randomisation and no ports



rand bit [1:0]in;

bit out;

//constraint wr_rd_en{wr_en != rd_en;};

endclass
