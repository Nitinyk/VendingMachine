class scoreboard;
	bit out;
endclass
